`timescale  1us/1us  //???? ???? ????
module xsfebpin_test;
  wire clk_out ;//????????,?????
  reg clk_in;// ???????,?????
  reg rst;
  xsfebpin u1(clk_in,rst,clk_out);//?????,???
  always #20 clk_in=~clk_in;
  initial
    begin
      clk_in=0;
      #100 rst=1;
      #200 rst=1;
      #400 rst=0;
      #6000 $stop;
    end
  initial $monitor($time, , ,"clk_in=%b  clk_out=%b",clk_in,clk_out);
endmodule
