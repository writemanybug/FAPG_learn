`timescale  1us/1us  //???? ???? ????
module div_3;
  wire out ;//????????,?????
  reg clk;// ???????,?????
  reg res;
  reg[7:0] n;
  jifenping u1(out,clk,res,n);//?????,???
  always #20 clk=~clk;
  initial
    begin
      clk=0;
      n=7;
      #100 res=1;
      #200 res=1;
      #400 res=0;
      #6000 $stop;
    end
  initial $monitor($time, , ,"clk=%b  out=%b",clk,out);
endmodule
