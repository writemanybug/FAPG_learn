library verilog;
use verilog.vl_types.all;
entity xsfebpin_test is
end xsfebpin_test;
