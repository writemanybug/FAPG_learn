library verilog;
use verilog.vl_types.all;
entity factor is
end factor;
