`timescale  1us/1us  //???? ???? ????
module counter_test;
  wire[4:0] out ;//????????,?????
  reg clk,rst;// ???????,?????
  counter u1(clk,rst,out);//?????,???
  always #20 clk=~clk;
  initial
    begin
      clk=0;rst=0;
      #50 rst=1;
      #6000 $stop;
    end
  initial $monitor($time, , ,"clk=%b rst=%b out=%b",clk,rst,out);
endmodule