library verilog;
use verilog.vl_types.all;
entity led_test is
end led_test;
