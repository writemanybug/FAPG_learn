library verilog;
use verilog.vl_types.all;
entity encoder8_3_test is
end encoder8_3_test;
