library verilog;
use verilog.vl_types.all;
entity stop_test is
end stop_test;
