library verilog;
use verilog.vl_types.all;
entity erfenpin_test is
end erfenpin_test;
