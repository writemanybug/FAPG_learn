library verilog;
use verilog.vl_types.all;
entity div_3 is
end div_3;
