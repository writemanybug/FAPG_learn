`timescale  1us/1us  //???? ???? ????
module erfenpin_test;
  wire out ;//????????,?????
  reg clk;// ???????,?????
  erfenpin u1(clk,out);//?????,???
  always #20 clk=~clk;
  initial
    begin
      clk=0;
      #6000 $stop;
    end
  initial $monitor($time, , ,"clk=%b  out=%b",clk,out);
endmodule
